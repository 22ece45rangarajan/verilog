module pipo_tb();
  reg [3:0]d;
  reg res,clk,load;
  wire [3:0]y;
  pipo  dut(d,res,clk,load,y);
  always #5 clk= ~clk;
  initial begin
    $monitor("time=%t,d=%b,res=%b,clk=%b,load=%b,y=%b",$time,d,res,clk,load,y);
  load=0;d=4'b0000;res=1;clk=0;
  #5;res=0;
  #10;d=4'b1001;load=1;
  #5;load=0;
  #15;d=4'b1010;load=1;
  #5;load=0;
  end
  initial begin
    $dumpfile("tvk.vcd");
    $dumpvars;
    #50 $finish;
  end
endmodule
