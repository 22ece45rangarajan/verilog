module encoder_8x3_tb();
  reg [7:0]a;
  wire [3:0]b;
  encoder_8x3 dut (a,b);
  initial begin
    $monitor("time=%0t,a=%b,b=%b",$time,a,b);
       a=8'b00000000;
    #5;a=8'b00011100;
    #5;a=8'b00001000;
    #5;a=8'b00010000;
    #5;a=8'b00100000;
    #5;a=8'b01000000;
    #5;a=8'b10000000;
  end
  initial begin
    $dumpfile("TVK.vcd");
    $dumpvars(0,encoder_8x3_tb);
    #50 $finish;
  end 
endmodule
