module dff(d,res,clk,q);
  input d,res,clk;
  output reg q;
  always @ (posedge clk)begin
    if (res)
      q<=0;
    else
      q<=d;
  end 
endmodule
